library ieee;
use ieee.std_logic_1164.all;

entity ejemplo1git is
	port(
			x1, x2: in std_logic_vector(3 downto 0);
			displays: out std_logic_vector(13 downto 0) 
			);
end ejemplo1git;
architecture bev of ejemplo1git

begin
--TODO
end bev;
