--cambio
library ieee;
use ieee.std_logic_1164.all;
entity adder is
	port(
			x1, x2 : in std_logic_vector(3 downto 0);
			result: out std_logic_vector(3 downto 0);
			carry : out std_logic_vector
			);
end adder;
architecture bev of adder

begin
--TODO
end bev;
